// must file (Do not delete)
